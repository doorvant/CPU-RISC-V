`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/07/13 11:38:14
// Design Name: 
// Module Name: RF
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module RF(
    input clk,
    input rst_n,
    input [4:0] rR1,
    input [4:0] rR2,
    input [4:0] wR_wb,
    input rf_we_wb,
    input [31:0] wD,
    output reg [31:0] rD1,
    output reg [31:0] rD2
    );
    
    reg [31:0] x0 = 32'h00000000;
    reg [31:0] x1 = 32'h00000000;
    reg [31:0] x2 = 32'h00000000;
    reg [31:0] x3 = 32'h00000000;
    reg [31:0] x4 = 32'h00000000;
    reg [31:0] x5 = 32'h00000000;
    reg [31:0] x6 = 32'h00000000;
    reg [31:0] x7 = 32'h00000000;
    reg [31:0] x8 = 32'h00000000;
    reg [31:0] x9 = 32'h00000000;
    reg [31:0] x10 = 32'h00000000;
    reg [31:0] x11 = 32'h00000000;
    reg [31:0] x12 = 32'h00000000;
    reg [31:0] x13 = 32'h00000000;
    reg [31:0] x14 = 32'h00000000;
    reg [31:0] x15 = 32'h00000000;
    reg [31:0] x16 = 32'h00000000;
    reg [31:0] x17 = 32'h00000000;
    reg [31:0] x18 = 32'h00000000;
    reg [31:0] x19 = 32'h00000000;
    reg [31:0] x20 = 32'h00000000;
    reg [31:0] x21 = 32'h00000000;
    reg [31:0] x22 = 32'h00000000;
    reg [31:0] x23 = 32'h00000000;
    reg [31:0] x24 = 32'h00000000;
    reg [31:0] x25 = 32'h00000000;
    reg [31:0] x26 = 32'h00000000;
    reg [31:0] x27 = 32'h00000000;
    reg [31:0] x28 = 32'h00000000;
    reg [31:0] x29 = 32'h00000000;
    reg [31:0] x30 = 32'h00000000;
    reg [31:0] x31 = 32'h00000000;
    
    always @(rR1) begin
            case(rR1)
                5'd00: rD1 = 32'h00000000;
                5'd01: rD1 = x1;
                5'd02: rD1 = x2;
                5'd03: rD1 = x3;
                5'd04: rD1 = x4;
                5'd05: rD1 = x5;
                5'd06: rD1 = x6;
                5'd07: rD1 = x7;
                5'd08: rD1 = x8;
                5'd09: rD1 = x9;
                5'd10: rD1 = x10;
                5'd11: rD1 = x11;
                5'd12: rD1 = x12;
                5'd13: rD1 = x13;
                5'd14: rD1 = x14;
                5'd15: rD1 = x15;
                5'd16: rD1 = x16;
                5'd17: rD1 = x17;
                5'd18: rD1 = x18;
                5'd19: rD1 = x19;
                5'd20: rD1 = x20;
                5'd21: rD1 = x21;
                5'd22: rD1 = x22;
                5'd23: rD1 = x23;
                5'd24: rD1 = x24;
                5'd25: rD1 = x25;
                5'd26: rD1 = x26;
                5'd27: rD1 = x27;
                5'd28: rD1 = x28;
                5'd29: rD1 = x29;
                5'd30: rD1 = x30;
                5'd31: rD1 = x31;
            endcase
    end
    
    always @(rR2) begin
            case(rR2)
                5'd00: rD2 = 32'h00000000;
                5'd01: rD2 = x1;
                5'd02: rD2 = x2;
                5'd03: rD2 = x3;
                5'd04: rD2 = x4;
                5'd05: rD2 = x5;
                5'd06: rD2 = x6;
                5'd07: rD2 = x7;
                5'd08: rD2 = x8;
                5'd09: rD2 = x9;
                5'd10: rD2 = x10;
                5'd11: rD2 = x11;
                5'd12: rD2 = x12;
                5'd13: rD2 = x13;
                5'd14: rD2 = x14;
                5'd15: rD2 = x15;
                5'd16: rD2 = x16;
                5'd17: rD2 = x17;
                5'd18: rD2 = x18;
                5'd19: rD2 = x19;
                5'd20: rD2 = x20;
                5'd21: rD2 = x21;
                5'd22: rD2 = x22;
                5'd23: rD2 = x23;
                5'd24: rD2 = x24;
                5'd25: rD2 = x25;
                5'd26: rD2 = x26;
                5'd27: rD2 = x27;
                5'd28: rD2 = x28;
                5'd29: rD2 = x29;
                5'd30: rD2 = x30;
                5'd31: rD2 = x31;
            endcase
    end

    always @(posedge clk or negedge rst_n) begin
        if(rst_n == 1'b0) begin
            x0 <= 32'h00000000; 
            x1 <= 32'h00000000; 
            x2 <= 32'h00000000; 
            x3 <= 32'h00000000; 
            x4 <= 32'h00000000; 
            x5 <= 32'h00000000; 
            x6 <= 32'h00000000; 
            x7 <= 32'h00000000; 
            x8 <= 32'h00000000; 
            x9 <= 32'h00000000; 
            x10 <= 32'h00000000;
            x11 <= 32'h00000000;
            x12 <= 32'h00000000;
            x13 <= 32'h00000000;
            x14 <= 32'h00000000;
            x15 <= 32'h00000000;
            x16 <= 32'h00000000;
            x17 <= 32'h00000000;
            x18 <= 32'h00000000;
            x19 <= 32'h00000000;
            x20 <= 32'h00000000;
            x21 <= 32'h00000000;
            x22 <= 32'h00000000;
            x23 <= 32'h00000000;
            x24 <= 32'h00000000;
            x25 <= 32'h00000000;
            x26 <= 32'h00000000;
            x27 <= 32'h00000000;
            x28 <= 32'h00000000;
            x29 <= 32'h00000000;
            x30 <= 32'h00000000;
            x31 <= 32'h00000000;
        end           
        else if(rf_we_wb == 1'b1)
            case(wR_wb)
                5'd00: x0 <= 32'h00000000;
                5'd01: x1 <= wD;
                5'd02: x2 <= wD;
                5'd03: x3 <= wD;
                5'd04: x4 <= wD;
                5'd05: x5 <= wD;
                5'd06: x6 <= wD;
                5'd07: x7 <= wD;
                5'd08: x8 <= wD;
                5'd09: x9 <= wD;
                5'd10: x10 <= wD;
                5'd11: x11 <= wD;
                5'd12: x12 <= wD;
                5'd13: x13 <= wD;
                5'd14: x14 <= wD;
                5'd15: x15 <= wD;
                5'd16: x16 <= wD;
                5'd17: x17 <= wD;
                5'd18: x18 <= wD;
                5'd19: x19 <= wD;
                5'd20: x20 <= wD;
                5'd21: x21 <= wD;
                5'd22: x22 <= wD;
                5'd23: x23 <= wD;
                5'd24: x24 <= wD;
                5'd25: x25 <= wD;
                5'd26: x26 <= wD;
                5'd27: x27 <= wD;
                5'd28: x28 <= wD;
                5'd29: x29 <= wD;
                5'd30: x30 <= wD;
                5'd31: x31 <= wD;
            endcase    
    end  
    
endmodule
